           A     A     A     A     A     A     A     A     A     A     A     A     A_    A_    A     A     A     A     A     A     A     A_    A     A     A     A     A     A     A     A_    A_    A_    A_    A_    A_    A_    A_    A     A     A/    A     A/    A_    A_    A_    A_    A_    A_    A(    A_    A)    A_    A_    A_    A_    A     !A/    !A     !A_    !A_    !A_    !A/    !A     !A_    !A     !A\    !A/    !A     !A_    !A_    !A/    !A     !A_    !A_    !A_    !A/    !A     !A/    !A     !A_    !A_    !A_    !A/    !A/    'A     'A/    'A_    'A_    'A/    'A     'A     'A_    'A_    'A/    'A     'A/    'A_    'A/    'A     'A/    'A     'A     'A/    'A     'A(    'A_    'A_    'A     'A     'A)    'A     'A\    -A_    -A_    -A_    -A/    -A\    -A_    -A_    -A_    -A/    -A\    -A_    -A_    -A/    -A_    -A/    -A     -A     -A/    -A_    -A/    -A_    -A_    -A_    -A_    -A/    -A     -A     -A_    3A_    3AC    3A     3AT    3Ae    3At    3Ar    3Ai    3As    3A_    3A_    3A_    3A_    3A     3A_    3A_    3A_    3A     3A_    3A_    3A     3A_    3A     3A     3A     3A     3A     3A