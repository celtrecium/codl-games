         #A⣨  #A⢦  #A⣤  #A⢮  #A⡀  #A⠸  #A⠹  #A⣛  #A⢛  #A⡻  #A⠹  #A