
      ⣠  FA⣾  FA⣿  FA⣿  FA⣿  FA⣿  FA⣿  FA⣿  FA⣷  FA⣄  FA⣿  FA⣿  FA⣿  FA⣿  FA⠿  FA⠿  FA⣿  FA⣿  FA⣿  FA⣿  FA⣿  FA⣿  FA⣿  FA⠁  FA     FA   FA⠈  FA⣿  FA⣿  FA⣿  FA