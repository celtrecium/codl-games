P      *    A     A     A     A     A     A     A.    A     A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A,    A     A     A     A     A     A.    A     A     A     A     A     A     A     A     A,    A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A,    A     A     A     A.    A       .    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A,    A     A     A     A     A     A     A     A     A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A*    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A            A     A.    A     A     A     A     A     A     A     A     A.    A     A     A     A     A     A     A     A*    A     A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A*    A     A     A     A     A     A     A     A     A     A*    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A,    A            A     A     A     A     A     A*    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A*    A     A     A     A     A     A     A     A     A     A     A     A*    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A,    A     A     A     A     A     A     A     A.    A     A     A     A     A     A     A     A     A.    A     A     A     A.    A     A            A     A     A     A     A     A     A     A     A     A.    A     A     A     A     A,    A     A     A     A.    A     A     A     A     A     A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A     A     A.    A     A     A     A     A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A,    A     A     A     A     A     A     A     A            A*    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A,    A     A     A     A     A     A     A*    A     A     A     A     A     A     A     A     A     A     A*    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A.    A            A     A     A     A     A*    A     A     A     A     A     A     A     A     A     A     A     A     Ao    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A*    A     A     A     A     A,    A     A     A     A     A     A     A     A     A,    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A            A     A     A     A     A     A     A     A     A     A     A     A     A     A*    A     A     A     A     A     A     A     A.    A     A     A     A     A*    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A*    A     A     A     A     A     A     A     A     A     A     A     A     A     Ao    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A.    A     A     A     A     A            A,    A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A,    A     A     A     A.    A     A     A*    A     A     A     A     A     A     A     A     A     A     A     A*    A     A     A     A     A*    A     A     A     A     A     A     A     A     A     A     A*    A     A     A     A     A     A     A     A     A*    A     A     A     A            A     A     A     A     A     A     A     A*    A     A     A     Ao    A     A     A,    A     A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A.    A     A     A     A,    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A,    A     A     A     A     A     A     A       *    A     A     A     A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A,    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A,    A     A     A     A.    A     A     A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A     A     A.    A            A     A     A     A     A     A     A     A     A     A.    A     A     A     A     A     A     A     A     A     A,    A     A     A     A     A     A     A.    A     A     A     A,    A     A     A     A     A     A     A.    A     A     A     A     A.    A     A     A     A     A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     Ao    A     A     A.    A     A     A     A     A     A            A     A     A     A     A     A     A     A     A     A     A     A     A     A*    A     A     A     A     A     A     A     A.    A     A     A     A     A*    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A*    A     A     A     A     A     A     A     A     A     A     A     A     A     Ao    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A            A.    A     A     A     A     A     A,    A     A     A     A     A     A     A     A     A     A     A     A*    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A*    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A.    A     A     A     A     A     A     A     A     A            A     A     A     A     A     A     A     A     A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     Ao    A     A     A     A     A     A,    A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A,    A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A.    A            A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A.    A     A.    A     A     A     A     A     A     A     A     A     A     A     A     A,    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A*    A     A     A     A     A*    A     A     A     A     A     A     A     A     A     A     A*    A     A     A     A     A     A     A     A     A*    A     A     A     A     A            A     A     A     A     A     A     A     A     A     A     A.    A     A     A     A     A     A     A     A*    A     A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A*    A     A.    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A.    A     A     A     A     A     A     A     A,    A            A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     Ao    A     A     A     A     A     A     A     A     A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A,    A     A     A     A     A     A     A     A     A,    A     A     A     A     A     A     A     A     A     A     A     A     A            A     A     A.    A     A*    A     A     A     A     A     A     A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A,    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A*    A     A     A     A     A     A     A     A     A     A,    A     A     A     A     A     A            A     A     A     A     A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A     A,    A     A     A     A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A.    A     A     A     A     A.    A     A     A     A     A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     Ao    A     A     A     A     A     A     A.    A     A            A,    A     A     A     A     A     A     A     A     A     A     A     A     A     A,    A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A,    A     A     A     A     A     A     A     A     A     A     A     A            A     A     A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A,    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A.    A     A     A     A     A.    A     A     A     A     A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A       *    A     A     A     A     A     A     A.    A     A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A,    A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A,    A     A     A     A     A            A     A     A     A     A     A     A*    A     A     A     A     A     A     A     A     A     A     A     A     A*    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A*    A     A     A     A     A     A     A     A     A     A     A     A     A     Ao    A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A     A,    A            A,    A     A     A,    A     A     A     A     A     A.    A     A     A     A     A,    A     A     A     A     A     A     A     A     A     A     A     A     A.    A     A     A     A     A     A     A     A     A     A     A.    A     A     A     A     A     A     A     A     A     A.    A     A     A.    A     A     A     A     A     A     A     A.    A     A     A     A     A     A     A,    A     A     A     A,    A     A     A     A     A.    A     A     A       