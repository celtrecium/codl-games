      /    #A~    #A~    #A~    #A\    #A     #A\    #A-    #AV    #A-    #A/    #A       