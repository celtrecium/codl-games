      /    &A_    &A_    &A_    &A\    &A            &A/    &A     &A\    &A              