
           FA.    FA-    FA-    FA-    FA-    FA-    FA-    FA.    FA       |    FA     FA     FA_    FA_    FA_    FA_    FA     FA     FA|    FA|    FA_    FA'    FA     FA     FA     FA     FA'    FA_    FA|    FA